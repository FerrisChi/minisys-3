`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

module Idecode32 (
	input			reset,
    input			clock,
    output	[31:0]	read_data_1,	// ����ĵ�һ������
    output	[31:0]	read_data_2,	// ����ĵڶ�������
    input	[31:0]	Instruction,	// ȡָ��Ԫ����ָ��
    input	[31:0]	read_data,		// ��DATA RAM or I/O portȡ��������
    input	[31:0]	ALU_result,		// ��ִ�е�Ԫ��������Ľ������Ҫ��չ��������32λ
    input			Jal,			// ���Կ��Ƶ�Ԫ��˵����JALָ�� 
    input			RegWrite,		// ���Կ��Ƶ�Ԫ
    input			MemtoReg,		// ���Կ��Ƶ�Ԫ
    input			RegDst,			// ���Կ��Ƶ�Ԫ
    output	[31:0]	Sign_extend,	// ���뵥Ԫ�������չ���32λ������
    input	[31:0]	opcplus4		// ����ȡָ��Ԫ��JAL����
);
    
    reg[31:0] register[0:31];			   //�Ĵ����鹲32��32λ�Ĵ���
    reg[4:0] write_register_address;        // Ҫд�ļĴ����ĺ�
    reg[31:0] write_data;                   // Ҫд�Ĵ��������ݷ�����

    wire[4:0] read_register_1_address;    // Ҫ���ĵ�һ���Ĵ����ĺţ�rs��
    wire[4:0] read_register_2_address;     // Ҫ���ĵڶ����Ĵ����ĺţ�rt��
    wire[4:0] write_register_address_1;   // r-formָ��Ҫд�ļĴ����ĺţ�rd��
    wire[4:0] write_register_address_0;    // i-formָ��Ҫд�ļĴ����ĺ�(rt)
    wire[15:0] Instruction_immediate_value;  // ָ���е�������
    wire[5:0] opcode;                       // ָ����
    
    assign opcode = Instruction[31:26];	//OP
    assign read_register_1_address = ������//rs 
    assign read_register_2_address = ������//rt 
    assign write_register_address_1 = ������// rd(r-form)
    assign write_register_address_0 = ������//rt(i-form)
    assign Instruction_immediate_value = ������//data,rladr(i-form)


    wire sign;                                            // ȡ����λ��ֵ

    assign sign = ������
    assign Sign_extend[31:0] = ������
    
    assign read_data_1 = ������
    assign read_data_2 = ������
    
    always @* begin                                            //�������ָ����ָͬ���µ�Ŀ��Ĵ���

    end
    
    always @* begin  //������̻�������ʵ�ֽṹͼ�����µĶ�·ѡ����,׼��Ҫд������
 
     end
    
    integer i;
    always @(posedge clock) begin       // ������дĿ��Ĵ���
        if(reset==1) begin              // ��ʼ���Ĵ�����
            for(i=0;i<32;i=i+1) register[i] <= 0;
        end else if(RegWrite==1) begin  // ע��Ĵ���0�����0


        end
    end
endmodule
